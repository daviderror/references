`timescale 1ns / 1ps

module heart_beat_tb;

    initial begin
        $stop();
    end
endmodule
